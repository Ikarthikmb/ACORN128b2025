module ch_fn(
	input x, y, z,
	output ch_out
);
	// LAB Problem-1: Correct ch_out here
	assign ch_out = 'b0;
	
endmodule
